//
//
//

package pkg_classes;


// include for all classes implementation
  
`include "transaction.sv"
`include "output_transaction.sv"
`include "Stimulus.sv"
`include "input_monitor.sv"
`include "output_monitor.sv"
`include "GoldModel.sv"
`include "Checker"
//`include "Coverage.sv"
`include "tb_overall.sv"
`include "interface.sv"
endpackage


