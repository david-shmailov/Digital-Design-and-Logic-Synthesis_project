Module Decoder (
            input   rst,
                    clk,
                    DATA_IN,

            output  data_out,


            );


            
endmodule